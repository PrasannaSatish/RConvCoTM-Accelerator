module axi_gpio_o_1 (
    // AXI clock & reset 
    input s_axi_aclk,
    input s_axi_aresetn,

    // GPIO output 
    output [0:0] gpio_io_o
);

endmodule