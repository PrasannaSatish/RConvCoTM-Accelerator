
// AXI-Stream Interface Skeleton (Data Path Only)

module axis_if #
(
    parameter DATA_WIDTH = 32
)
(
    input  wire                     clk,
    input  wire                     rst_n,

    input  wire                     ACLK,
    input  wire                     ARESETN,

    // AXI-Stream Slave Interface (Input to Accelerator)
    input  wire [DATA_WIDTH-1:0]    S_AXIS_TDATA,
    input  wire                     S_AXIS_TVALID,
    output wire                     S_AXIS_TREADY,
    input  wire                     S_AXIS_TLAST,

    // AXI-Stream Master Interface (Output from Accelerator)
    output wire [DATA_WIDTH-1:0]    M_AXIS_TDATA,
    output wire                     M_AXIS_TVALID,
    input  wire                     M_AXIS_TREADY,
    output wire                     M_AXIS_TLAST
);

  

endmodule
