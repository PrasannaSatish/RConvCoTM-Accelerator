module dma 
(
	input m_tready,
	output [127:0] m_tdata,
	output [15:0] m_tkeep,
	output m_tlast,
	output m_tvalid 
);

endmodule
