`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 14.07.2025 13:02:46
// Design Name: 
// Module Name: class_top_tb
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////

module class_top_tb;
    reg clk;
    reg rst;
    reg [18:0]model_params;
    reg [14:0]count = 0;
    reg [127:0] total_img;
    wire [31:0]bram_addr_a;
    wire [31:0]bram_addr_a2;
    wire tready;
    reg tvalid;
    reg [15:0]tkeep;
    reg tlast;
    reg [3:0]label;
    reg [3:0]calc_label;
    reg [255:0]clause_write;
    reg [255:0]weight_write;
    wire enb;
    wire [31:0]web ;
    wire [255:0] dinb;
    reg [20:0] success;
    reg [20:0] fail;
    reg opm;
    wire [3:0]output_params;
    
     initial clk = 0;
    always #5 clk = ~clk;
    integer img_count = 0;
    class_top
    uut
    (clk,rst,model_params,total_img,clause_write,weight_write,tvalid,tkeep,tlast,bram_addr_a,bram_addr_a2,tready,enb,output_params,web,dinb);
    initial 
    begin    
        count = 0;
        success = 0;
        fail = 0; 
        tvalid = 1;
        rst = 1;
        model_params = 19'b1010_010001100_001_101;
        #100
        rst = 0;
        #10
//number 0
       #10 total_img = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
       #10 total_img = 128'b00000000000000000000000000000000011110000111000000000000000000001111111110000000000000000000111111100000000000000000011100000000;
       #10 total_img = 128'b00000111000001110000000000000001110000001110000000000000001110000001110000000000000001100000011100000000000000001111000111000000;
       #10 total_img = 128'b00000000011000000001100000000000000011000000001100000000000000011000000001100000000000000011000000001100000000000000011000000000;
       #10 total_img = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000110000000000000000110000000110;
       #10 total_img = 128'b00000000000000000000000000000000000000000000000000000000001111101111000000000000000011100001110000000000000000111000000011000000;
       #10 total_img = 128'b00000000000000000000000000000000000000000000000000001111111000000000000000000000000111111110000000000000000000000000000000000000;
       #10 total_img = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
end
        always @(posedge clk) begin
        if (tready)begin
       if(count == 0)begin
       count <= count + 1; 
        total_img = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
       end
       if(count == 1)begin
       count <= count + 1; 
       total_img = 128'b00000000000000000000000000000000011110000111000000000000000000001111111110000000000000000000111111100000000000000000011100000000;
       end
       if(count == 2)begin
       count <= count + 1; 
       total_img = 128'b00000111000001110000000000000001110000001110000000000000001110000001110000000000000001100000011100000000000000001111000111000000;
       end
       if(count == 3)begin
       count <= count + 1; 
       total_img = 128'b00000000011000000001100000000000000011000000001100000000000000011000000001100000000000000011000000001100000000000000011000000000;
       end
       if(count == 4)begin
       count <= count + 1; 
       total_img = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000110000000000000000110000000110;
       end
       if(count == 5)begin
       count <= count + 1; 
       total_img = 128'b00000000000000000000000000000000000000000000000000000000001111101111000000000000000011100001110000000000000000111000000011000000;
       end
       if(count == 6)begin
       count <= count + 1; 
       total_img = 128'b00000000000000000000000000000000000000000000000000001111111000000000000000000000000111111110000000000000000000000000000000000000;
       end
       if(count == 7)begin
       count <= count + 1; 
       total_img = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
       end
        if(count == 8)begin
       count <= count + 1; 
        total_img = 128'b00000000000000000000000000000000000000000000000000001111111000000000000000000000000111111110000000000000000000000000000000000000;
       end
       if(count == 9)begin
       count <= count + 1; 
       total_img = 128'b00000000000000000000000000000000011110000111000000000000000000001111111110000000000000000000111111100000000000000000011100000000;
       end
       if(count == 10)begin
       count <= count + 1; 
       total_img = 128'b00000111000001110000000000000001110000001110000000000000001110000001110000000000000001100000011100000000000000001111000111000000;
       end
       if(count == 11)begin
       count <= count + 1; 
       total_img = 128'b00000000011000000001100000000000000011000000001100000000000000011000000001100000000000000011000000001100000000000000011000000000;
       end
       if(count == 12)begin
       count <= count + 1; 
       total_img = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000110000000000000000110000000110;
       end
       if(count == 13)begin
       count <= count + 1; 
       total_img = 128'b00000000000000000000000000000000000000000000000000000000001111101111000000000000000011100001110000000000000000111000000011000000;
       end
       if(count == 14)begin
       count <= count + 1; 
       total_img = 128'b00000000000000000000000000000000000000000000000000001111111000000000000000000000000111111110000000000000000000000000000000000000;
       end
       if(count == 15)begin
       count <= count + 1; 
       total_img = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
       end
       
       
       end
       end
       always @(posedge clk) begin
          case (bram_addr_a)
        
            0: clause_write = 142'b0010001100000000000000000000000000000000000000010000100001000001000001000000000000000100001000000000000010001011100000001100010000001000000000;
            1: clause_write = 142'b0011100000000000000000001000000000000000000000000000000000000000000100000000000011000000000001000000000001001001000001111100001000010000100000;
            2: clause_write = 142'b0000000000000000000000010110111110000000000000000000100000000000000000100001100110111111011111000000000000000000101110000000000000000100011000;
            3: clause_write = 142'b1100000000000000000000001100000000000000000000000000000000000000000011000001111101110111011011000000001101011111111111111101111111111111100000;
            4: clause_write = 142'b1111111111000000000000011111111111100000000000001111111110111011100110000000000000000111111101000000000000011111111110000000000000000000000000;
            5: clause_write = 142'b0000000000000000000000000000000000000000000000000000000001000100001000000000010100001000000000000000000000010100010100001100011000100001100011;
            6: clause_write = 142'b0000000000000000000000000000100000010001000000001000000000000000000000000000001100000000000010000000000000000000000000000000000000001001011001;
            7: clause_write = 142'b0111100000000000000000011111111100000000000000000000001101110011001100000000000111010110111111000000000000011001100100100010000100000000100010;
            8: clause_write = 142'b0000000000000000000001000000000000000000000000000010000000010000100000000000000000000000000000000000000001000000000000010000000000001000000000;
            9: clause_write = 142'b0111111011111111110100011010100000000000000000000000000000000000000000100000000000000000000001000000000000011111111001110111000010101110011100;
            10: clause_write = 142'b1111110111100000000000011101110011110011100000100001000010000000000000000000000000001101101111000000000000000000111110000100111001110111101111;
            11: clause_write = 142'b0000000000000000000000011111100000000000000000000000000000000000000000101111111111011111111111000000011101111111110111111111111010111111101000;
            12: clause_write = 142'b1000000000000000000000011111111100000000000000000000000000100111111111100011111111111111111111000000000000011111111111011111011000000000000000;
            13: clause_write = 142'b0011111111111111000000011111110000000000000000011100000000000000000000000000000000000000000111000000000011011111111100000000001101111101111011;
            14: clause_write = 142'b1111111111010000000000010100101100100000000000001000000100000000000000000000000000000001111011000000000000000001111110000010000101001111011110;
            15: clause_write = 142'b1100000000000000000000011110000000000000000000000000000000000000000000100011001111111111101101000001011110001010001111001100110111111111111110;
            16: clause_write = 142'b1110000000000000000000000110010000000000000000000000100001000100000000000000000110010010100000000000000000010000010000001100001000110001100110;
            17: clause_write = 142'b1111111111111000000000011111111111111111110000110001100011000100000000000000000000000001111111000000000000000000000110001100011001110011100111;
            18: clause_write = 142'b1101101110010101000111011111111001000000000000010000100001000000000000000000000000000000000001000000000000000010101110000000001000111111001101;
            19: clause_write = 142'b1111110111110011100000001111101111001011100000100000000000000000000000000000000000000000010111000000000000000000011110111101111111111011111111;
            20: clause_write = 142'b0000000000000000100000100000000000100000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            21: clause_write = 142'b1111111011111111000000011111001111101100000000000010001011000000000000000000000000000000000000000000000000000000011111100000000000000000101111;
            22: clause_write = 142'b0000001010000000000000000001101001010000000000010000000001000111110000000000000000000101000000000000000000000010000000000100011000000000000000;
            23: clause_write = 142'b1110110001111111110000010000000000000000000000000010000100001000000000000000000000000000000111000101010111101111011010000001000111001010011111;
            24: clause_write = 142'b1111110000000000000000011111111111111100000000100001000010000100001000000000000111111111111111000000000000000011111110011100111001110011100111;
            25: clause_write = 142'b1111011111111110000000011011111100000000000000000010001000001001110011000000000000000000011111000000000001111111111111100000000110001000010000;
            26: clause_write = 142'b1111111101111111111000000000000000000000000000000010000100000000000000000000000000000000000001001111111110111111101111110011100011101111001111;
            27: clause_write = 142'b1000000000000000000000011111111111111111100000000000000000000000001000000111111111111111101111000000000000000000111101111111111111111110100111;
            28: clause_write = 142'b0000000000000100000000000000000110000000000000110000011000000001000010000000000000000000000000000000000000000100000000000000000000001000000001;
            29: clause_write = 142'b1111100000000000000000011111111111111111100000000000000000000000000000000000111111111111111111000000000000000000111111111111111111111111111111;
            30: clause_write = 142'b0000001000000000000000000000010000000000000000000001000010000110010110000000000010000100100000000000000000001000000000000000100000000000000000;
            31: clause_write = 142'b0000000101010000110000000111001000000000000000100000000000000100000000000000000000000000000000000000000000101100011000001000001000100000100011;
            32: clause_write = 142'b1000000000000010100000000001000110000000000000100001000010000100000000100000000000000000000000000000000000010100000010000000000001000000000000;
            33: clause_write = 142'b0000000000000000000000000111110000000000000000000000000000001000010000100111001101011100100001000000000000011101111011111000100001000000011000;
            34: clause_write = 142'b0000000000100000000000000000000000010000000000000010000100000000000000000000000000010000000001000000000000000000000001000000000100001000011000;
            35: clause_write = 142'b1111111111100000000000000000000000000000000000000000000000000000000000100000000000000111111111001111111111111111111111111111111111101110011100;
            36: clause_write = 142'b1000000000000000000000011111111111111000000000000000000000000001111111100011111111111111111111000000000000000111111111111111111111110000000000;
            37: clause_write = 142'b1111111111111111111110011000000000000000000000000110000000000000000000000000000000000000000001000011111111111111111111100011100111111111111111;
            38: clause_write = 142'b0001000110110000000000000001001000000000010000100000100000100001000100000000000000000000101010000000000000000000000100000000000000010000000000;
            39: clause_write = 142'b1100000000000000000000011110000000000000000000000000000000000000010000100001111111111111111111000001111111111111111111111111111111111110011100;
            40: clause_write = 142'b1111000000000000000000000111111101010110000000000000000000000000001000000000111111101110101111000000000000000000001101111111011011111110101111;
            41: clause_write = 142'b1100000000000000000000000011011100000000000000000000000100000000000000000000011110101110100100000000000000001111011111100001000100000001000111;
            42: clause_write = 142'b0001000100000000000000010000000000000000000000011000000000000101110000100000000000100000000000000000000100000001000000000000001000000000000000;
            43: clause_write = 142'b1101010111010000000000000010000100110000000000000001000000000000000000000000000000000001011101000000000000001010101110000000011001100100011011;
            44: clause_write = 142'b1111111111111110000000011111111111111111100000000000000000000000000000000000000000000011111111000000000000000001111111111111111111111111111111;
            45: clause_write = 142'b1100000000000000000000011011111010100000000000000000000011011000000000100000111010100101111111000000000000000001101101111100000000000000010100;
            46: clause_write = 142'b0000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000100000000000000000000000000000000000000000000000;
            47: clause_write = 142'b0101010000000000000000010011000001000010000000000110000000000000000000000000000000010010000000000000000000000000000000000000000000001100000011;
            48: clause_write = 142'b0001000010101000000000000000000000000000000000100000000000000000000000000000000000000110010000000000000011010000000000001100000000010001100010;
            49: clause_write = 142'b1111000100100010000000010110000000000000000000000100001100011000010000000000000000000000000110000000101010110100110010100001000000001000001000;
            50: clause_write = 142'b1000001110011000000000001101010101001010100100000000000010000000000000000000000000000011100001000000000000000000000000000100000000000001011001;
            51: clause_write = 142'b1111111100000000000000011000000000000000000000000010000000000000000000000000000001111111111111000011111111111111111111110011100111001111111111;
            52: clause_write = 142'b1111111000000000000000011111111101111111111000100001000010000100001000000000000001111111111111000000000000000000000010011100111001110011100111;
            53: clause_write = 142'b1000000000000000000000010000000000000000000000000000000000000100001000000000000000000000011000000000000011010101111111111100001000110000100011;
            54: clause_write = 142'b1111101110100110000000010101110100000000000000000110110011000000011000100000000000000000101011000000000000000111111000000000000000000000000000;
            55: clause_write = 142'b1111111000000000000000011011111111010110110000000001000010000000000000000000000011111101011111000000000000000000000110111100111010110011101111;
            56: clause_write = 142'b1000000000000000100000000000000000000000000000000000000000000000000010000000000000000000000000000000000100000000000001000011110000011000000000;
            57: clause_write = 142'b1111010101101000000000000110100000000000000000011000100010000100001000000000000000000001110100000000000001111010110100000000000000000011000011;
            58: clause_write = 142'b0000000000000000000000000000000000001000000000000000000100000000000000000000001000000000000000000000000000000000000000110010000010000000010000;
            59: clause_write = 142'b1111111111111111111100011000000000000000000000000010000100001000000000000000000000000000000010000001111111111111111111100011100111101111111111;
            60: clause_write = 142'b1111000000000000000000011111111111011000000000110000110001100011100011000000000011111011111101000000000000000011111110001100001000010000000000;
            61: clause_write = 142'b0000000000000000000000000000000000000000000000000000000000010000000000001000000000000000000000000000000000000000000000000000000000000000000000;
            62: clause_write = 142'b1111111111111111111100011111110000000000000000111110011100000000000000000000000000000000000001000000000111111111111110000000000111111111111011;
            63: clause_write = 142'b1111111111111111110000011000000000000000000000000010000000000000000000000000000000000000000111000111111111101111111111110011110111111111111111;
            64: clause_write = 142'b1110110000000000000000010110001011110001110000110000000010000000000000000000000011010101010101000000000000000000000110000000011000110111110011;
            65: clause_write = 142'b0000000001000011100000000010000000000010000000001000000000000000000000000000000000000000000000000000000000000000000000000010000100000110100111;
            66: clause_write = 142'b0111111111100110101010001111110000000000000000000011000010000000000000000000000000000000000000000000000001110111011010000000000000011111001111;
            67: clause_write = 142'b1011100000000000000000010011101110000100000000000000000000000000000000100000000011101111001011000000000000000000001010111101101001100100000000;
            68: clause_write = 142'b0000000000000001000001000000101100000000000000000000000100100000000000000000000000000000000000000000000000000000000000010000000000000000000000;
            69: clause_write = 142'b1111111111111111111000011111111000000000000000111111110000000000000000000000000000000000000011000000000001111111111110000000000000111111111111;
            70: clause_write = 142'b0111111100000000000000011100000000000000000000000000000000010000100011000000000000111111010110000001111111111011111111110001100110001000010000;
            71: clause_write = 142'b0100000000000000000000011111111000000000000000000000000000000011001111100011101111111111101111000000000001011111111111111111110111010000000000;
            72: clause_write = 142'b0001000011000000000000001001000100000000000000000110000100000000000000000000000000000011110000000000000010000110000001100000000100001000011000;
            73: clause_write = 142'b1111111111110000000000011111111111111110000000110000100001100011000110000000000000000011111111000000000000000001111110000100001000010000100001;
            74: clause_write = 142'b0011100000000000000000000011010111000000000000000000000000000000001011100000000101000001010000000000000000000000000001000010101010010000000000;
            75: clause_write = 142'b1000110001101000000000000000001101100000000000000000100001100000000010000000000000000000010001000000000000001111000100001000001000110000000000;
            76: clause_write = 142'b1100000000000000000000011111100000000000000000000000000000000000000000100111111111111111111111000000001111111111111111110111111111111111111110;
            77: clause_write = 142'b1111110111100000000000011000000000000000000000000010000100011000100001100000000000001111111111000001101110101110011111010011000101000100010000;
            78: clause_write = 142'b1101011111111000000000011011110000000000000000000000000000000000010001100000000000000111001101000000000001111111111111111111110111001000010000;
            79: clause_write = 142'b0000000000000000000000000000000000000000000000000000100000000000001000000000000000000000000100000000010000000000000000000000000000000010000000;
            80: clause_write = 142'b1011111111101011011101011110011100000000000000011010000000000000000000000000000000000000000000000000000001110111111111000001000111111011111011;
            81: clause_write = 142'b0000000000000000000000000000000000000000000000000010010000000000000000000000000110010010100000000000000110001000000100000010000100001000111111;
            82: clause_write = 142'b0000000000000000000000011100000000000000000000000000000000000000000000100111111111111111111111000001111111111111111111111111111111111111011100;
            83: clause_write = 142'b0101011011111011101111000001000000000000000000100000000010000100000000000000000000000000000000000000000000000000011000001100011000110000000011;
            84: clause_write = 142'b0000000100010000000000000000000101000000000000000000000000000000000000000000000000000100110000000000000000000100001000101110101010011000000001;
            85: clause_write = 142'b1101110000000000000000000110001001110000000000011100101011010010101100000000000000010110111110000000000000000111110100000000000000000000100001;
            86: clause_write = 142'b1100000000000000000000011111110000000000000000000000000000011011111100000001111111111111111111000000000111111111111111111111110000000000000000;
            87: clause_write = 142'b0100000000000000000000001000100000000000000000000000000000001000001000000001100010001111010001000000000000101111010010000000000000000000000111;
            88: clause_write = 142'b1000011001000000000000001001000000000000000000000010011101100000000111000000000000011101100110000000000111011010011001100000000000000000000000;
            89: clause_write = 142'b1111111111110111000000011101111110000000000000100001000110000100001001100000000000000000000010000000000000000111111110000000000000000000000000;
            90: clause_write = 142'b0111100000000000000000011011111111011111010110000001100000000000000000000000000000010111100100000000000000000000000000000000011000010000000010;
            91: clause_write = 142'b1101000000000000000000000101111101101000000000100111110100001000110011000000000000101111011110000000000000000000011100000000000000001000010000;
            92: clause_write = 142'b0000000010000000000000000000000000010000000000000000000000000010000010000000000000000100000000000000000000000100000001100000100000100000100000;
            93: clause_write = 142'b1010000000000000000000011110111101010000000000000000000000110101111111100001111010011011110110000000000000000001111111110110101000000000000000;
            94: clause_write = 142'b1111111111111111111000011111111111110000000000000010001001110110000000000000000000000000000001000000000000000011111111100000000000000000100111;
            95: clause_write = 142'b1101001000001001100000000111101010000000000000110100001100001000000000000000000000000000000111000000000000000000001000000000000000001010011011;
            96: clause_write = 142'b1111111111111111111000011111111100000000000000000000000000000000000000000000000000000000000111000000000011111111111111111111111111111111111111;
            97: clause_write = 142'b0100000000000000000000000000011011000000000000000000000000000110000010000000010100100100010011000000000000011100010000000001001001100000100001;
            98: clause_write = 142'b1110101111010101111000010001101111111111101100100000000000000000000000000000000000000000000010000000000000000000000000011111111111111011111111;
            99: clause_write = 142'b1111110000000000000000011111111111111100000000000000000000000000000000000000000111111111111111000000000000000001111111111111111111111111111111;
            100: clause_write = 142'b1111111111111111110000011111011111111110000000110001100000000000000000000000000000000000000111000000000000000001111110001100011011110111111111;
            101: clause_write = 142'b0000000000000000000000000000000001001000000000110010000000000000000000000000000011000000000000000000000000000000000000000000000000001100000011;
            102: clause_write = 142'b0000010100101000000000000000000000000000000000000000000000000000000100000000000000000001100000000000000011000000010000000001111100010000100000;
            103: clause_write = 142'b1111100000000000000000011111111111011111111110000000000000000000001000000000000111111111111111000000000000000000000001111100111001110011100111;
            104: clause_write = 142'b0001000000000000000000000000000000000001000000000000000000000000010000000000000000100000000000000000000000000000000001000000000100000000001000;
            105: clause_write = 142'b0001000000000000000000000000000000000000000000000000000000000000001000000000001000000000100000000000000100001000000000000000011000000001000000;
            106: clause_write = 142'b0111110101111000000000011111000000000000000000000000000000000000000001100000000000000001111110000000010111101011111110111110010011111110010000;
            107: clause_write = 142'b0000000000000000000000000000000000000010000000000010000000000000000000000000000000000000000000000000000000000000000000000001000000001010000110;
            108: clause_write = 142'b1001010000000000000000001000010000000000000000000000000001000011000001100000000001011000000010000000000000101001000000000000000000100000010000;
            109: clause_write = 142'b1000000000000000000000011111111111111110000000000000000000000000001000000111111111111111111111000000000000000011111111111111111111111111100111;
            110: clause_write = 142'b1110111111111111100000011011111111011000000000000110001100111111100110000000000000000000001111000000000000000000011110100000000000000000000000;
            111: clause_write = 142'b1111111111000000000000001110000000000000000000000000000000000000000011000000000000000111111110000000011111110111111110111111101111001100000000;
            112: clause_write = 142'b1000000000000000000000010010000101000000000100000000000000000010000000000000100010011001100000000000000000000000000000100100010100010000000000;
            113: clause_write = 142'b1100000000000000000000011111111110000000000000000000000000000000000011100011111111111111111111000000000000111111111111111111111111111111011000;
            114: clause_write = 142'b1010110110100000000000010111101111100000000000001101100100001000000000000000000000001111111110000000000000000111101110000000000000001100001000;
            115: clause_write = 142'b1111111001010101110111111110010010011110000000100000000000000000000000000000000000000000000000000000000000000001011100110101111101011111010110;
            116: clause_write = 142'b0000000010000000000000000000000000001000000000000000010000000000000000000000000000001000000000000000000000000000001000000000001001101000000000;
            117: clause_write = 142'b1111111111111111100000011111110000000000000000000000000000000000000000000000000000000000111111000000011111111111111111111111111111111111111111;
            118: clause_write = 142'b0000000010001100000000000000000000000000000000000000000000000001000000000000000000000000000000000000010000000000000001011000001000010000000000;
            119: clause_write = 142'b0100101110000000000000010111101000000000000000000100001000100001000010000000000000010100111010000000000011011000100110100011000100000000100000;
            120: clause_write = 142'b0000000000000000000000000000000110111000000000010000000000000000000000000000111000000110100001000000000000000000000110000100000000010001011101;
            121: clause_write = 142'b1111111101100000000000011000000000000000000000000100001000010000110000100000000000000011111111000000110011111111111111100011000111000110011100;
            122: clause_write = 142'b0000000111100000000000000010000001101010000000000000100000000000000000000000000000000000000000000000000000000000000000110100000000011011111010;
            123: clause_write = 142'b0001000000000001001000000001010001100000000000000000000100000000000000000000000000000000000001000000000000000000000000010000000110001010000010;
            124: clause_write = 142'b0000000000000000000000000010000000000000000000100000000010000010000010100000000000001010000010000000001000000000001010000000011000000000000000;
            125: clause_write = 142'b0101010100100000000000010010000101111100000000001100000010000000000000000000000000001111001011000000000000000000000001000000000000000011100000;
            126: clause_write = 142'b0110000000000000000000001100000000000000000000000000000000110001110001100000101100100010010011000000000000111110111101111010001100001000010000;
            127: clause_write = 142'b0000000000000000000000000000000000000000000000000000000001000000000100000000000100000100001001000000000001100000000000001000010000000001000011;
            128: clause_write = 142'b0001001110011000000000011111111000000000000000000110011001100110001000000000000000000010100101000000000011111111011000000010000000000000000000;
            129: clause_write = 142'b0001110110000011110000000000000000000000000000000000000000000000000001000000000000000000000000000000000011000100100001000000000001111000010000;
            130: clause_write = 142'b1001000010010011000000000000100111100000000000100001000000000100000001100000000000000000000110000000000000000000010100000000010000000000000000;
            131: clause_write = 142'b1000000000000000000000010011111111111000000000000000000000000000010001000000011110011111111111000000000000000000011011111101010111001100011000;
            132: clause_write = 142'b0000000000000000000000000000000000000000000100000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            133: clause_write = 142'b1110000000000000000000000011101101110000000000000000000011000000000000000000000011011111010111000000000000000000000001111100001000010000111111;
            134: clause_write = 142'b0000000010100000000000000000001000000000000000000000010000011000000000000000000000000101011000000000000010000000000000000010000100000100001111;
            135: clause_write = 142'b1111111111111111110000011111000000000000000000000010000000000000000000000000000000000000000111000000011111111111101111110011110111111111111111;
            136: clause_write = 142'b0111110111100000000000011110111111111111000000000100001000100011001100000000000000001111001110000000000000000000001010000000000000000000100000;
            137: clause_write = 142'b0000000000000000000000000000000000000000000000011000000100001000001100000000000100000001100000000000000000000000000000000000000010000000000000;
            138: clause_write = 142'b1111100000000000000000010111000000000000000000000000000000000000010011100000011111101111111111000000001111111111111111110111111111101110011000;
            139: clause_write = 142'b1111111111111111111111011111111111111111000000110000000000000000000000000000000000000000000000000000000000000000111110001100111111111111111111;
        
          endcase
        end
        
        always @(posedge clk) begin
  case (bram_addr_a2)

    0: weight_write = 256'b0000000000000000100100000111100000000000101101110100000000100000000001010001010101111011101000000000000000000000001111110010110100100000000000001110000001000100000000001110100000100011001110001010111000001101101101011100011100111100011111000000000000000000;
    1: weight_write = 256'b0000000000101010111010101111101010111001011101100110011110110100000000000101010100100001001011010000000000000001101000000101000011010100000000010000000000000000000111011011001000100000000000000110100000000100000000000000000111111010100000000001001101110000;
    2: weight_write = 256'b0000000000001100110101000000000000000000000000001000000000000000001000000000000000000000000000010111000100110100000000111111011110000000000000000000100010000100110010111011111000011011110000110000000000110001100000000000010001000011110101110010100000000001;
    3: weight_write = 256'b0000000000000000000000000100000000001011110100000000100000000000000000000000000000000000010001001000000000011110110000000000001010101000000100011000001000000000000000000101100111000000000000111010000001111011110111000000000000000000000000000000000000100000;
    4: weight_write = 256'b0000000000000000000011101111100000010011101011010000000000101101100001000111110110011000001100111011000000000001100011000000000000000000010101111000010011000000000010000000000000000000000000001111111100011001010000000000000110100000000000000000011011101100;
    5: weight_write = 256'b0000000000000100000000000000011000000000000000000010001101100000000100000000010010011000000000010001110000000000100111100000000000010011010000010100000000000110001100100000000111111101100000000000000000000011011000000000000000000000000000000000000000000000;
    6: weight_write = 256'b1000010001001001101011101010000000000000000000000000010000000000000000000000111010000000010000000001010101000000000000000101000101001100000000000110110000000000000000000011010100000000000011000011000000000100000000011111001010000000000000000010000000000000;
    7: weight_write = 256'b0000000000001000000001000000000000000000000000000110000010000000000000000000000000000000000001000000001000000001011000111000000000000000000000000000000000000010110100000000000000000001000000000000000000000000000000000001100100111000000001000000000000000000;
    8: weight_write = 256'b0000000000000000100000000001100111100000000001011101100000000000000000000000000000000000000000000000000000000000000000000000100000000000000100000000000000000000011011010000000000000000000101100110000001001000000000011100011000000000000000000000000000100000;
    9: weight_write = 256'b0000000000000000000011011001000000010000011110010000000000111110100010010110111101110000000000000000001110001100000000000000000000000000010000000011001011100000000000111101100000000000000000000000000011001000010000000010000000000000000000000000001110111100;
    10: weight_write = 256'b1100000011100111000010000000011011101010001100011100000000001011101100000000110000010000000000011010101000000000110000000011010101100000000111101010100000000100000000110010111000011011001110001000000000010011011000000000000010111100000000000011100011110000;
    11: weight_write = 256'b0000000011100000101000111001101001100011011111101100000010010100000000011100010111010001101001000001110001101010010100000101011110011000000000010100001000000000000001110000111101100000000011111111011111111010000000000000000110000000000000000001000000101001;
    12: weight_write = 256'b1100000000001000000001000111110000000000000000000011001110000000000101011000000000000000000000011101001110111100000100001000000000000011101101010110101101101110011001000000001111010101000101100000000000000000000111000111111100010001101000101101100000000001;
    13: weight_write = 256'b0000000000000000100001111111101110101101010100000000100110100000000000000000000000000000001111101000000000000000000000000000100000000111110101100000000011010110111100100000001011000000000111101001000000011000000000000000000011010101000000000000000000010100;
    14: weight_write = 256'b0000000000000000000010000000011111101100011010100111011111111000011100100011111010101011000000010001100000000001100011000000000001111100110000000000000110100000000000001011000000000001101111000000000010000000001110011011110100000000000010000000010000000000;
    15: weight_write = 256'b0100000000000011000000000110010000000000100000000010001101001101000100000000100000000000000000000000000000000000100010000100000000100000000111110101100000000001100110001100001000101001110101100001010101100000000011001011100000000001110101000011100000000000;
    16: weight_write = 256'b0000000010000000001010111101011111000101100110000000000000000100000000001001000011010001101000101000111000111010001000000101010000000000000000011010111000000000000001110000100110100000000000000100011111101101101110100000000111111010100000000011110011101101;
    17: weight_write = 256'b0000000000000100000110010011010000000000000000001000000000000000001000000000101010100000000000001000010010011010000101100010101000000000001101010110101101101000000001000000001011111011011111100000000000000000000000000001110000100011010100010100010000000001;
    18: weight_write = 256'b0000000000000000100000000111101001010001011101101000111111111000000000000000000000000000011010010000000000111110010000000000000000000111101011100000000010010001100000000111100100000000000000101010111011101101000011011100011000000000000000000000000000100000;
    19: weight_write = 256'b0000000000000000000010000000011111111011010010101001000100010011111100100011010100100110001010000000000000000000000000000000000010000000001001101100000001000000000000101000100000000000000000000000000000011100010000000000101000001111111100000000000000000000;
    20: weight_write = 256'b0000010011100000100100100001000010111000100011000100000000000101100001100010110111000010001110000000000000000000000011100100000000010101000000000010010110110000101001111101000110001111000010100001010101111010110001100001100000000001010111011110001010001110;
    21: weight_write = 256'b0111011000010111000000000010000000000110001010000000000100000100000000010000000000001100100000000000000000000101111000000101010111001000000000000101011100000000010000000010010011100000000000000110100000000110000000000000000100010100000000000000001101110000;
    22: weight_write = 256'b0000000000000010001110001101000000000000000000000100011110000000001000000000000000000000000000000110001000000001101110000000000010110000100111011011000000000011111101111101011101111000100000100000000000111100010000000000000010011000000001000000000000000000;
    23: weight_write = 256'b0000000000000000010100100110010001100000000010000010001101100000000000000000000000000000000000000000000000000000000011110001011100100000000100101100001101111100100000000100000000000000000110101010111111101100000000000000000000000000000000000000000000100000;
    24: weight_write = 256'b0000000000000000000000101000000000010011111110000101101110000000000000100011100111010000000010000000000000000001100011000000000000000000000011110011101000001111111110111101000000000000110001100000000000100100010000000000101000000000000001111110010000000000;
    25: weight_write = 256'b0100011010010000100100000100011000000000010011010000011011001101000000010110111001110000000000010001110000000000000001001000000000100000000111111111111110011000001000000111000111110110001011110001010101101100000001101111000000000000011101000011100000000000;
    26: weight_write = 256'b0000000010000000000000000000110000101000000000010100111101111100000000010000000011010001100000010000000000010110011100000011110111111100000000011000100100000000001010111000001110000000000000000101000000000101101100100000000111110100100000000010001101001001;
    27: weight_write = 256'b0000000000000011110110001011010000000000000000000000000000000000000011010010000000000000000000000101000011101100000111100001010001000000010000000001101010111000000001101010110010010011100100010000000000000000000011100010000100010011010101000000000000000001;
    28: weight_write = 256'b0000000000000000100000000000010101001010001100000000000100111000000000000000000000000000111011111000000000111110010000000000001010101000000001010001000010011111111110011010111100000000000000110101000001001100000000000000000000000000000000000000000000100000;
    29: weight_write = 256'b0000000000000000000011100111111111101110000000000100001110101101100000000100101101100100111110010110000000000000000000000000000011101010101000011100000110100000000000011001100000000000000000000000000000011001010000000010101110100000000000000000000000000000;
    30: weight_write = 256'b0000000000000000000000001001011000000000010011010000000000100000000010000111001111111001011110000000000000000000001000110100000000011000001000010111100000000100000000001010011111100110111000001000000000100000000000000000000000000000011101000000000000000000;
    31: weight_write = 256'b0000000010000000000000000000000000000101100100001100100110100000000000010000000001001011000011100111100011100111100100000101000111001100000000001011100100000000010000000010000000000000000011111111000000000110010110000000000100101001000000000001000000110000;
    32: weight_write = 256'b0110000000001000000001000000000000000000000000001000000000111110110110110010000000000000000000011001100001011011111110011000000000000000001101010111000000001110011000000000001000000001110000110000000000000000000110001100001011010000101111001000010000000001;
    33: weight_write = 256'b0000000000000000001010010000110110100000000100000000001101000011111111000000000000000000100000000000000000100000000011000110000000000000000100111110100000000000100000000010101001000000000000110010000001111110111001000000000000000000000000000000000000010110;
    34: weight_write = 256'b0000000000000000000000010110111111010000010100110000000010101101100001011111110001100000000000000000000000000000000000000000000010000000010000000000010100100000000010000000000000000001011111100000000010000000000101110110000000000000000000000000010000000000;
    35: weight_write = 256'b1101100011101100000000000010010000000000100000000011000100000011000100000000100000000000000000000000000000000000111010011000000000000000000110101011000000000001001001111010001110101111110100000000000000001000111001101111010001011100000000000000000000000000;
    36: weight_write = 256'b0111111000111001111110100000000000010110110011101100010111110000000000000111000011101000000000000000000000011010001011001101000000000000000000011000100100000000010000000000100011001110001100000110100000000100000000000000000110111110000000000011011100011001;
    37: weight_write = 256'b0000000000001111111011000000000000000000000000000100111010001110011000000000000000000000000001011001111000000000001000010010001010000011101101010110000000001110000001101010110100111010100111000000000000000000000000000001000000001000000000101101100000000000;
    38: weight_write = 256'b0000000000000000100111111000011101010001011010001000100000000000000000000000000000000000000000000000000000000000000000000000111000000000000100111110100000000000110010110000000000011111111111010001110111111000000000000000000011101100000000000000000000100000;
    39: weight_write = 256'b0000000000000000000000001010000000010000010100100001000111001101111100100011100001010000000011000111100000000000000000000000000000000000000011110000000100100000000010000000000000000000000000000000000011101011110000000001000000100000000000000000010000000000;
    40: weight_write = 256'b0000010011100001101111110000110000000000000110001100000000111110111001011010100110111000000000000000000000000000101100001100000000100010110000001110010011111001001001111010001000010010001000111010111000100000000000000000100000000001010111000000000000000000;
    41: weight_write = 256'b0101011110011011010000000010000000010000000010000000000011001001111111100111011100011011011110110100000000010000000000000101011100011100000000010000000000000000000111001100100101000000000000000110100000000100000000000000000111100101100000000010000000000000;
    42: weight_write = 256'b0110000000000001000000100011000000000000000000000000000000000000001000000000000000000000000001100111100101001000000010100011011110000000000000000000001110011000000000000000001110001111100100010000000000000000000000000000010001110010001101000000000000000000;
    43: weight_write = 256'b0000000000000000010001110110110100000011111111010101010001101000000000000000000000000000001001000000000000000000000000000000101001101000000100000001011101111100001011110001110100000000000000110010000001111000000000000000000000000000000000000000000000010110;
    44: weight_write = 256'b0000000000000000000000010010000000010000001110100010010001001010100000101101000100000100111101101011101110001100000000000000000000000000010000000011111111000000000001001011000000000010000000000000000000101101011100111011011011000000000010000000000100111000;
    45: weight_write = 256'b0000000000000100000000110000110001010101111111101101001001000100000010100000100000000000000000010001110000000000001010010100000000000000000000010001001101100010001111110010111000100110100000000000000000000101000000000100100000000001111000000000000001011110;
    46: weight_write = 256'b1000001000010010010000000000000000010011011011101100011101011100000000010000000100001000000000000000000000010100001111111101100001101100000000011011110100000000011110010010111100001110001100000110100000000100000000000000000101010100000000000010000000010000;
    47: weight_write = 256'b0010000000000010101010101000100000000000000000001000000000000000000000000000111101100000000001000000001000000000001000110010111000110110001101010110000000000000110011101010110100101010001101100000000000000000000000000000001000011000000001000000000000000000;
    48: weight_write = 256'b1111111000000000010101001000101000000001000010001000001010011000000000000000000000000000000000000000000000000000000000000000000000000000000100110111001100000000101011110100000000000000000110001110000001111100000000000000000000000000000000000000000000100010;
    49: weight_write = 256'b0000000000000000000000111110100000010000001110111100001010000000000001110110111101100110001010000000000000000000000000000000000000000000001010101011111010100000000000010000100000000010000000000000000000100001110000000000011000000000000000000000010000000001;

  endcase
end

//        always @(posedge output_params[4]) begin
//        count = count + 1;
//        #10
//        prst[1] = 1'b1;
//        #10 prst[1] = 1'b0;
//        #10
//             if(count == 1)begin
////         //number 1
//         total_img = 512'b00000000000000000000011000000000000000000000000001100000000000000000000000000111000000000000000000000000011000000000000000000000000011100000000000000000000000001110000000000000000000000000111000000000000000000000000011100000000000000000000000001110000000000000000000000000111000000000000000000000000011100000000000000000000000001110000000000000000000000000011000000000000000000000000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
//        #10
//           total_img = 512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000000000000000000000000111000000000000000000000000011100000000000000000000000000111000000000000000000000000011100000000000000000000000001110000;     
//        end
//        else if(count == 2)begin
//         //number 2
//         total_img = 512'b10000000000000000000011111000000000000000000000011110000000000000000000000011111000000000000000000000011111000000000000000000000001111000000000000000000000001111000000000000000000000000111000000000000000000000000011100000000000000000000000011100000000000000000000000000110000000000000000000000000011000000000000000000000000001100000000000000000000000000111000000000000000000000000001111010000000000000000000000011111100000000000000000000000011100000000000000000000000000000000000000000000000000000000000000000000;
//        #10
//           total_img = 512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000011110000000000000111111111111111000000000000111111111111111100000000000001000000111111;     
//        end
//        else if(count == 3)begin
//         //number 3
//         total_img = 512'b00000000000000000110000000000000000000000000011100000000000000000000000000111100000000000000000000000001111100000000000000000000000011100000000000000000000000011100000000000000000000000001100000000000000000000000001100000000000000000000000000100000000000000000000000000110000000110000000000000000011000000111000000000000000001100001111000000000000000000111111111000000000000000000001111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
//        #10
//           total_img = 512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111100000000000000000000111111111000000000000000000011100011100000000000000000011000000110000000000000000001100000110000000000000000000110000010000;     
//        end
//        else if(count == 4)begin
//         //number 4
//         total_img = 512'b11000000000000000111111111111100000000000000011100000111100000000000000000110000111100000000000000000011100011100000000000000000001110011110000000000000000000110011110000000000000000000011001110000000000000000000001101110000000000000000000000111110000000000000000000000011111000000000000000000000011111000000000000000000000001111100000000000000000000000111100000000000000000000000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
//        #10
//           total_img = 512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100000000000000000000000000111000000000000000000000000011100000000000000000000000001110000000000000000000000000111111111111000000000000000011111111111;     
//        end
//        else if(count == 5)begin
//         //number 5
//         total_img = 512'b10000000000000001100000000011000000000000000110000000001000000000000000011100000000000000000000000000111100000000000000000000000001111111110000000000000000000001111111000000000000000000000000001100000000000000000000000000110000000000000000000000000111000000000000000000000000011000000000000000000000000011100000000000000000010001111100000000000000001111111111100000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
//        #10
//         total_img = 512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111000000000000000000011111111110000000000000000011110000111100000000000000001110000000110000000000000001110000000011000000000000000110000000001;     
//        end
//        else if(count == 6)begin
//         //number 6
//         total_img = 512'b00000000000000111110111111110000000000000011101111111111000000000000001111111110111100000000000000111111100011110000000000000011111100001111000000000000000000000001111000000000000000000000000111100000000000000000000000111100000000000000000000000111110000000000000000000001111110000000000000000000100111110000000000000000000111111110000000000000000000111111110000000000000000000011111100000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
//        #10
//           total_img = 512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111000000000000000000001111111110000000000000000011111111111100000000000000011111111111110000000000000001111101111111;     
//        end
//        else if(count == 7)begin
//         //number 7
//         total_img = 512'b00000000000000000011100000000000000000000000011100000000000000000000000001110000000000000000000000000110000000000000000000000000111000000000000000000000000011000000000000000000000000011100000000000000000000000001110000000000000000000000000110000000001111000000000000011111111111111111100000000000111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
//        #10
//           total_img = 512'b00000000000000000000000000000000000000001110000000000000000000000001111000000000000000000000000001100000000000000000000000001110000000000000000000000000111000000000000000000000000011100000000000000000000000011100000000000000000000000001110000000000000000000000001110000000;     
//        end
//        else if(count == 8)begin
//         //number 8
//         total_img = 512'b00000000000000000000111111100000000000000000000011111100000000000000000000001111100000000000000000000001111110000000000000000000001111111000000000000000000001111111100000000000000000001111001110000000000000000001111000011100000000000000000111000111110000000000000000111111111110000000000000000011111111110000000000000000001110000000000000000000000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
//        #10
//           total_img = 512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000000000000000000000001111110000000000000000000001111111000000000000000000001111011100000000000000000001111001110000000000000000000111000110000000000000000000011101111;     
//        end
//        else if(count == 9)begin
//         //number 9
//         total_img = 512'b00000000000000000011100000000000000000000000001110011111000000000000000000110011111100000000000000000111011111111000000000000000011111100011100000000000000001111000001100000000000000001111000001110000000000000000111000011110000000000000000111100111110000000000000000011111111100000000000000000000111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
//        #10
//           total_img = 512'b00000000000000000000000000000000000000000001110000000000000000000000001111000000000000000000000001111000000000000000000000000111000000000000000000000000011000000000000000000000000011100000000000000000000000001100000000000000000000000001110000000000000000000000000111000000;     
////        end
//always @(posedge opm) begin
//    label = (img_count)/96;
//    if(label == calc_label)success = success + 1;
//    else fail = fail + 1;
//    #10 prst[1] = 1'b1;
//    #10 prst[1] = 1'b0;
//    #10 load_next_chunk();
//    #10 load_next_chunk();
//end
//always @(posedge clk) begin
//calc_label = output_params[3:0];
//opm <= output_params[4];
//end
//reg [511:0] total_img;
//integer fd, r;
//reg [1024*8:1] line; // buffer for each line
//reg [783:0] bits784;
//integer j;
//integer cycle_count = 0;

//initial begin
//    fd = $fopen("1000testset.hex","r");
//    if (fd == 0) begin
//        $display("Error: could not open file");
//        $finish;
//    end
//end

//task load_next_chunk;
//        begin
//            if (cycle_count == 0) begin
//                // read one image = 784 ASCII chars
//                for (j=0; j<784; j=j+1) begin
//                    r = $fgetc(fd);
//                    if (r == "0")
//                        bits784[783-j] = 1'b0;
//                    else if (r == "1")
//                        bits784[783-j] = 1'b1;
//                    else
//                        j = j - 1; // skip newline or junk
//                end
//                // chunk 1 = lower 512
//                total_img = bits784[511:0];
//                cycle_count = 1;
//            end
//            else begin
//                // chunk 2 = upper 271 + padding
//                total_img = {241'b0, bits784[783:512]};
//                cycle_count = 0;
//                img_count = img_count + 1;
//            end
//        end
//    endtask
        
endmodule
